�� sr *com.win.tools.easy.common.PersitentManager�ۓ�~��  xr java.util.HashMap���`� F 
loadFactorI 	thresholdxp?@     w      t *com.win.tools.easy.platform.PlatFormConfigsr *com.win.tools.easy.platform.PlatFormConfigHC�F�Y I stateL disablePluginst Ljava/util/List;L frameBoundst Ljava/awt/Rectangle;xp    psr java.awt.Rectangleðj�jt I heightI widthI xI yxp  �    Q   �x